"000000000000000000000000000000000000000000" when "00000000",
"100000000000000000000000000000000000100001" when "00000001",
"000000000000000000000000000000000000000001" when "00000010",
"100000000000000000000000000000000000100010" when "00000011",
"000000000000000000000000000000000000000010" when "00000100",
"100000000000000000000000000000000000100011" when "00000101",
"000000000000000000000000000000000000000011" when "00000110",
"100000000000000000000000000000000000100100" when "00000111",
"000000000000000000000000000000000000000100" when "00001000",
"100000000000000000000000000000000010000000" when "00010001",
"000000000000000000000000000000000000000000" when "00010010",
"100000000000000000000000000000000010000010" when "00010011",
"000000000000000000000000000000000000000010" when "00010100",
"100000000000000000000000000000000010000011" when "00010101",
"000000000000000000000000000000000000000011" when "00010110",
"100000000000000000000000000000000010000100" when "00010111",
"000000000000000000000000000000000000000100" when "00011000",
"100000000000000000000000000000001000000000" when "00100001",
"000000000000000000000000000000000000000000" when "00100010",
"100000000000000000000000000000001000000001" when "00100011",
"000000000000000000000000000000000000000001" when "00100100",
"100000000000000000000000000000001000000011" when "00100101",
"000000000000000000000000000000000000000011" when "00100110",
"100000000000000000000000000000001000000100" when "00100111",
"000000000000000000000000000000000000000100" when "00101000",
"100000000000000000000000000000100000000000" when "00110001",
"000000000000000000000000000000000000000000" when "00110010",
"100000000000000000000000000000100000000001" when "00110011",
"000000000000000000000000000000000000000001" when "00110100",
"100000000000000000000000000000100000000010" when "00110101",
"000000000000000000000000000000000000000010" when "00110110",
"100000000000000000000000000000100000000100" when "00110111",
"000000000000000000000000000000000000000100" when "00111000",
"100000000000000000000000000010000000000000" when "01000001",
"000000000000000000000000000000000000000000" when "01000010",
"100000000000000000000000000010000000000001" when "01000011",
"000000000000000000000000000000000000000001" when "01000100",
"100000000000000000000000000010000000000010" when "01000101",
"000000000000000000000000000000000000000010" when "01000110",
"100000000000000000000000000010000000000011" when "01000111",
"000000000000000000000000000000000000000011" when "01001000",
"100000000000000000000000000000001010000000" when "00111001",
"000000000000000000000000000000000000000000" when "01000000",
"100000000010000000000000000000000000001000" when "01001001",
"000000000000000000000000000000000000001000" when "01001010",
"100000000000000010000000000000000000000000" when "00001001",
"000000000000000000000000000001000000000000" when "00011001",
"000000000000000000000000000100000000000000" when "00101001",
"100000000000000000000000000000000000001000" when "01100000",
"100000000000000000000000001000000000001000" when "01100001",
"000000000000000000000000000000000000001000" when "01100010",
"100000000000000000000000000000000000001001" when "01110000",
"100000000000000000000000001000000000001001" when "01110001",
"000000000000000000000000000000000000001001" when "01110010",
"100000000000000000000000000000000000001010" when "10000000",
"100000000000000000000000001000000000001010" when "10000001",
"000000000000000000000000000000000000001010" when "10000010",
"100000000000000000000000000000000000001011" when "10010000",
"100000000000000000000000001000000000001011" when "10010001",
"000000000000000000000000000000000000001011" when "10010010",
"100000000000000000000000000000000000001100" when "10100000",
"100000000000000000000000001000000000001100" when "10100001",
"000000000000000000000000000000000000001100" when "10100010",
"100000000000000000000000000000000000001101" when "01100011",
"100000000000000000000000000000000000001101" when "01100100",
"100000000000000000000000000000000000101101" when "01100101",
"000000000000000000000000000000000000001101" when "01100110",
"100000000000000000000000000000000000001101" when "01110011",
"100000000000000000000000000000000000001101" when "01110100",
"100000000000000000000000000000000010001101" when "01110101",
"000000000000000000000000000000000000001101" when "01110110",
"100000000000000000000000000000000000001101" when "10000011",
"100000000000000000000000000000000000001101" when "10000100",
"100000000000000000000000000000001000001101" when "10000101",
"000000000000000000000000000000000000001101" when "10000110",
"100000000000000000000000000000000000001101" when "10010011",
"100000000000000000000000000000000000001101" when "10010100",
"100000000000000000000000000000100000001101" when "10010101",
"000000000000000000000000000000000000001101" when "10010110",
"100000000000000000000000000000000000001101" when "10100011",
"100000000000000000000000000000000000001101" when "10100100",
"100000000000000000000000000010000000001101" when "10100101",
"000000000000000000000000000000000000001101" when "10100110",
"100000000100000000000000000000000000000101" when "01100111",
"100000000000000000000000000000000000000101" when "01101000",
"100000000000000000000000000000000000000101" when "01101001",
"100000000000000000000000000000000000100101" when "01101010",
"000000000000000000000000000000000000000101" when "01101011",
"100000000100000000000000000000000000000101" when "01110111",
"100000000000000000000000000000000000000101" when "01111000",
"100000000000000000000000000000000000000101" when "01111001",
"100000000000000000000000000000000010000101" when "01111010",
"000000000000000000000000000000000000000101" when "01111011",
"100000000100000000000000000000000000000101" when "10000111",
"100000000000000000000000000000000000000101" when "10001000",
"100000000000000000000000000000000000000101" when "10001001",
"100000000000000000000000000000001000000101" when "10001010",
"000000000000000000000000000000000000000101" when "10001011",
"100000000100000000000000000000000000000101" when "10010111",
"100000000000000000000000000000000000000101" when "10011000",
"100000000000000000000000000000000000000101" when "10011001",
"100000000000000000000000000000100000000101" when "10011010",
"000000000000000000000000000000000000000101" when "10011011",
"100000000100000000000000000000000000000101" when "10100111",
"100000000000000000000000000000000000000101" when "10101000",
"100000000000000000000000000000000000000101" when "10101001",
"100000000000000000000000000010000000000101" when "10101010",
"000000000000000000000000000000000000000101" when "10101011",
"100000000000000000000000000000000000010000" when "10110000",
"100000000000000000000000001000000000010000" when "10110001",
"100000000000000100000000000000000000010000" when "10110010",
"000000000000000000000000000000000000010000" when "10110011",
"100000000000000000000000000000000000010001" when "11000000",
"100000000000000000000000001000000000010001" when "11000001",
"100000000000000100000000000000000000010001" when "11000010",
"000000000000000000000000000000000000010001" when "11000011",
"100000000000000000000000000000000000010010" when "11010000",
"100000000000000000000000001000000000010010" when "11010001",
"100000000000000100000000000000000000010010" when "11010010",
"000000000000000000000000000000000000010010" when "11010011",
"100000000000000000000000000000000000010011" when "11100000",
"100000000000000000000000001000000000010011" when "11100001",
"100000000000000100000000000000000000010011" when "11100010",
"000000000000000000000000000000000000010011" when "11100011",
"100000000000000000000000000000000000010100" when "11110000",
"100000000000000000000000001000000000010100" when "11110001",
"100000000000000100000000000000000000010100" when "11110010",
"000000000000000000000000000000000000010100" when "11110011",
"100000000000001000000000000000000000010101" when "10110101",
"100000000000000000000000000000000000010101" when "10110110",
"100000000000000000000000000000000000010101" when "10110111",
"100000000000000000000000000000000000110101" when "10111000",
"000000000000000000000000000000000000010101" when "10111001",
"100000000000001000000000000000000000010101" when "11000101",
"100000000000000000000000000000000000010101" when "11000110",
"100000000000000000000000000000000000010101" when "11000111",
"100000000000000000000000000000000010010101" when "11001000",
"000000000000000000000000000000000000010101" when "11001001",
"100000000000001000000000000000000000010101" when "11010101",
"100000000000000000000000000000000000010101" when "11010110",
"100000000000000000000000000000000000010101" when "11010111",
"100000000000000000000000000000001000010101" when "11011000",
"000000000000000000000000000000000000010101" when "11011001",
"100000000000001000000000000000000000010101" when "11100101",
"100000000000000000000000000000000000010101" when "11100110",
"100000000000000000000000000000000000010101" when "11100111",
"100000000000000000000000000000100000010101" when "11101000",
"000000000000000000000000000000000000010101" when "11101001",
"100000000000001000000000000000000000010101" when "11110101",
"100000000000000000000000000000000000010101" when "11110110",
"100000000000000000000000000000000000010101" when "11110111",
"100000000000000000000000000010000000010101" when "11111000",
"000000000000000000000000000000000000010101" when "11111001",
"100000000000000000000000010000000001000000" when "00001100",
"000000000000000000000000000000000000000000" when "00001101",
"100000000000010000000000010000000001000000" when "00011100",
"000000000000010000000000000000000000000000" when "00011101",
"100000000000100000000000010000000001000000" when "00101100",
"000000000000100000000000000000000000000000" when "00101101",
"100000000000110000000000010000000001000000" when "00111100",
"000000000000110000000000000000000000000000" when "00111101",
"100000000001000000000000010000000001000000" when "01001100",
"000000000001000000000000000000000000000000" when "01001101",
"100000000001010000000000010000000001000000" when "01011100",
"000000000001010000000000000000000000000000" when "01011101",
"100000000001100000000000010000000001000000" when "01101100",
"000000000001100000000000000000000000000000" when "01101101",
"100000000001110000000000010000000001000000" when "01111100",
"000000000001110000000000000000000000000000" when "01111101",
"000000000000000001000000000000000000000000" when "10001110",
"000000000000000000100000000000000000000000" when "10101110",
"000000000000000000010000000000000000000000" when "11001110",
"000000000000000000001000000000000000000000" when "11101110",
"000000000000000000000100000000000000000000" when "10011110",
"000000000000000000000010000000000000000000" when "10111110",
"000000000000000000000001000000000000000000" when "11011110",
"000000000000000000000000100000000000000000" when "11111110",
"001000000000000000000000000000000000000000" when "00001110",
"010000000000000000000000000000000000000000" when "00011110",
"000010000000000000000000000000000000000000" when "00101110",
"000100000000000000000000000000000000000000" when "00111110",
"000000100000000000000000000000000000000000" when "01001110",
"000001000000000000000000000000000000000000" when "01011110",
"000000001000000000000000000000000000000000" when "01101110",
"000000010000000000000000000000000000000000" when "01111110",
