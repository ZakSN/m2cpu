library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity byte_to_text is port
(
	byte_in : in std_logic_vector(7 downto 0);
	line_out : out std_logic_vector(9 downto 0);
	line_sel : in std_logic_vector(4 downto 0)
);
end entity byte_to_text;

architecture a0 of byte_to_text is
	constant non_printing : integer := 32;
	constant char_set_size : integer := 112;
	signal lo : std_logic_vector(9 downto 0);
	type font_rom_array is array (0 to (char_set_size * 25) - 1) of std_logic_vector(9 downto 0);
	signal font_rom : font_rom_array;
	signal byte_num : integer;
	signal line_num : integer;
	signal c_t_p : integer;
	signal char_to_print : integer;

begin

	byte_num <= to_integer(unsigned(byte_in));
	line_num <= to_integer(unsigned(line_sel));
	-- assuming that all chars we recieve print as either a space or map to a printing char
	-- non printing chars (zero-width) need to be filtered out earlier. 
	-- by the time we get here we have to print something
	-- the next line ensures we print something predictable
	char_to_print <= (byte_num - non_printing) when (byte_num >= non_printing) AND (byte_num < (char_set_size + non_printing - 1)) else 0;
	line_out <= font_rom((char_to_print * 25) + line_num);
	
-- prototype char:
-- top five lines and bottom five lines are blanked for
-- text seperation
-- texh chars have a one pixel buffer on each edge (look at examples below)
--	"0000000000",
--	"0000000000",
--	"0000000000",
--	"0000000000",
--	"0000000000",
--	
--	"0000000000",
--	"0000000000",
--	"0000000000",
--	"0000000000",
--	"0000000000",
--	"0000000000",
--	"0000000000",
--	"0000000000",
--	"0000000000",
--	"0000000000",
--	"0000000000",
--	"0000000000",
--	"0000000000",
--	"0000000000",
--	"0000000000",
--	
--	"0000000000",
--	"0000000000",
--	"0000000000",
--	"0000000000",
--	"0000000000",


-- literal miles of font rom:
-- char are surrounded by "--{X" and "--X}"
-- where X is the particular char

	font_rom <=(
		--{SPACE
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--SPACE}
		--{!
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000000000",
		"0000000000",
		"0000110000",
		"0000110000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--!}
		--{"
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0111001110",
		"0111001110",
		"0110001100",
		"0110001100",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--"}
		--{#
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0011001100",
		"0011001100",
		"0011001100",
		"0011001100",
		"0111111110",
		"0111111110",
		"0011001100",
		"0011001100",
		"0011001100",
		"0111111110",
		"0111111110",
		"0011001100",
		"0011001100",
		"0011001100",
		"0011001100",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--#}
		--{$
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000110000",
		"0000110000",
		"0011111100",
		"0011111100",
		"0110110110",
		"0110110110",
		"0110110000",
		"0011111100",
		"0000110110",
		"0110110110",
		"0110110110",
		"0011111100",
		"0011111100",
		"0000110000",
		"0000110000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--$}
		--{%
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"1111110011",
		"1100110011",
		"1111110011",
		"0000001100",
		"0000001100",
		"0000001100",
		"0000110000",
		"0000110000",
		"0000110000",
		"0011000000",
		"0011000000",
		"0011000000",
		"1100111111",
		"1100110011",
		"1100111111",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--%}
		--{&
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0011111100",
		"0111111110",
		"0110000110",
		"0111000110",
		"0011111100",
		"0001111000",
		"0011110000",
		"0110110000",
		"0110110000",
		"0110011000",
		"0110011000",
		"0110011110",
		"0011111110",
		"0001110110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--&}
		--{'
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0001111000",
		"0001111000",
		"0000110000",
		"0000110000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--'}
		--{(
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000110",
		"0000001100",
		"0000110000",
		"0001100000",
		"0011000000",
		"0011000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0011000000",
		"0011000000",
		"0001100000",
		"0000110000",
		"0000001100",
		"0000000110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--(}
		--{)
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0110000000",
		"0011000000",
		"0000110000",
		"0000011000",
		"0000001100",
		"0000001100",
		"0000000110",
		"0000000110",
		"0000000110",
		"0000001100",
		"0000001100",
		"0000011000",
		"0000110000",
		"0011000000",
		"0110000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--)}
		--{*
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000110000",
		"0000110000",
		"0111111110",
		"0111111110",
		"0001111000",
		"0011001100",
		"0011001100",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--*}
		--{+
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0111111111",
		"0111111111",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--+}
		--{,
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000011110",
		"0000011110",
		"0000011000",
		"0000011000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--,}
		--{-
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0111111110",
		"0111111110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		---}
		--.{
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000110000",
		"0001111000",
		"0001111000",
		"0000110000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--.}
		--{/
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000011",
		"0000000011",
		"0000000011",
		"0000001100",
		"0000001100",
		"0000001100",
		"0000110000",
		"0000110000",
		"0000110000",
		"0011000000",
		"0011000000",
		"0011000000",
		"1100000000",
		"1100000000",
		"1100000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--/}
		--{0
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0011111100",
		"0111111110",
		"0110000110",
		"0110000110",
		"0110011110",
		"0110011110",
		"0110110110",
		"0110110110",
		"0110110110",
		"0111100110",
		"0111100110",
		"0110000110",
		"0110000110",
		"0111111110",
		"0011111100",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--0}
		--{1
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000110000",
		"0000110000",
		"0011110000",
		"0011110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0111111110",
		"0111111110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--1}
		--{2
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0011111100",
		"0011111100",
		"0110000110",
		"0110000110",
		"0000000110",
		"0000001100",
		"0000001100",
		"0000110000",
		"0000110000",
		"0011000000",
		"0011000000",
		"0110000000",
		"0110000000",
		"0111111110",
		"0111111110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--2}
		--{3
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0011111100",
		"0011111100",
		"0110000110",
		"0110000110",
		"0000000110",
		"0000000110",
		"0000001100",
		"0001111000",
		"0000001100",
		"0000000110",
		"0000000110",
		"0110000110",
		"0110000110",
		"0011111100",
		"0011111100",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--3}
		--{4
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000001100",
		"0000111100",
		"0000111100",
		"0011001100",
		"0011001100",
		"0011001100",
		"0110001100",
		"0110001100",
		"0110001100",
		"0111111110",
		"0111111110",
		"0000001100",
		"0000001100",
		"0000001100",
		"0000001100",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--4}
		--{5
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0111111110",
		"0111111110",
		"0110000000",
		"0110000000",
		"0110000000",
		"0011111000",
		"0011111000",
		"0000001100",
		"0000001100",
		"0000000110",
		"0000000110",
		"0000000110",
		"0000000110",
		"0111111100",
		"0111111100",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--5}
		--{6
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0011111100",
		"0011111100",
		"0110000110",
		"0110000110",
		"0110000000",
		"0110000000",
		"0110000000",
		"0111111100",
		"0111111100",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0011111100",
		"0011111100",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--6}
		--{7
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0111111110",
		"0111111110",
		"0000000110",
		"0000000110",
		"0000000110",
		"0000001100",
		"0000001100",
		"0000001100",
		"0000011000",
		"0000011000",
		"0000011000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--7}
		--{8
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0011111100",
		"0011111100",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0011111100",
		"0011111100",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0011111100",
		"0011111100",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--8}
		--{9
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0011111100",
		"0011111100",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0011111110",
		"0011111110",
		"0000000110",
		"0000000110",
		"0000000110",
		"0000000110",
		"0011111100",
		"0011111100",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--9}
		--{:
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000111000",
		"0000111000",
		"0000111000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000111000",
		"0000111000",
		"0000111000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--:}
		--{;
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000111000",
		"0000111000",
		"0000111000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000111000",
		"0000111000",
		"0000011000",
		"0000011000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--;}
		--{<
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000110",
		"0000001100",
		"0000011000",
		"0000110000",
		"0001100000",
		"0011000000",
		"0110000000",
		"1100000000",
		"0110000000",
		"0011000000",
		"0001100000",
		"0000110000",
		"0000011000",
		"0000001100",
		"0000000110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--<}
		--{=
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0111111110",
		"0111111110",
		"0000000000",
		"0000000000",
		"0111111110",
		"0111111110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--=}
		--{>
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0110000000",
		"0011000000",
		"0001100000",
		"0000110000",
		"0000011000",
		"0000001100",
		"0000000110",
		"0000000011",
		"0000000110",
		"0000001100",
		"0000011000",
		"0000110000",
		"0001100000",
		"0011000000",
		"0110000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		-->}
		--{?
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0011111100",
		"0011111100",
		"0110000110",
		"0110000110",
		"0000000110",
		"0000001100",
		"0000001100",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000110000",
		"0000110000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--?}
		--{@
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0111111110",
		"0111111110",
		"1100000011",
		"1100000011",
		"1100011111",
		"1100011111",
		"1100110011",
		"1100110011",
		"1100110011",
		"1100011111",
		"1100011111",
		"1100000000",
		"1100000011",
		"0111111110",
		"0111111110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--@}
		--{A
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000110000",
		"0001111000",
		"0011001100",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0111111110",
		"0111111110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--A}
		--{B
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0111111100",
		"0111111100",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110111100",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0111111100",
		"0111111100",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--B}
		--{C
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0011111100",
		"0011111100",
		"0110000110",
		"0110000110",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000110",
		"0110000110",
		"0011111100",
		"0011111100",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--C}
		--{D
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0111111100",
		"0111111100",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0111111100",
		"0111111100",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--D}
		--{E
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0111111110",
		"0111111110",
		"0110000000",
		"0110000000",
		"0110000000",
		"0111111110",
		"0111111110",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0111111110",
		"0111111110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--E}
		--{F
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0111111110",
		"0111111110",
		"0110000000",
		"0110000000",
		"0110000000",
		"0111111110",
		"0111111110",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--F}
		--{G
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0011111100",
		"0011111100",
		"0110000110",
		"0110000110",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110011110",
		"0110011110",
		"0110000110",
		"0110000110",
		"0011111100",
		"0011111100",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--G}
		--{H
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0111111110",
		"0111111110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--H}
		--{I
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0111111110",
		"0111111110",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0111111110",
		"0111111110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--I}
		--{J
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0111111110",
		"0111111110",
		"0000000110",
		"0000000110",
		"0000000110",
		"0000000110",
		"0000000110",
		"0000000110",
		"0000000110",
		"0000000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0011111100",
		"0011111100",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--J}
		--{K
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110001100",
		"0110001100",
		"0110001100",
		"0110011000",
		"0111110000",
		"0110011000",
		"0110001100",
		"0110001100",
		"0110001100",
		"0110000110",
		"0110000110",
		"0110000110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--K}
		--{L
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0111111110",
		"0111111110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--L}
		--{M
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0110000110",
		"0111001110",
		"0111001110",
		"0110110110",
		"0110110110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--M}
		--{N
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0110000110",
		"0111000110",
		"0111000110",
		"0110110110",
		"0110110110",
		"0110001110",
		"0110001110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--N}
		--{O
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0011111100",
		"0011111100",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0011111100",
		"0011111100",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--O}
		--{P
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0111111100",
		"0111111100",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0111111100",
		"0111111100",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--P}
		--{Q
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0011111100",
		"0011111100",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110110110",
		"0110110110",
		"0110011110",
		"0110001110",
		"0011111110",
		"0011111110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--Q}
		--{R
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0111111100",
		"0111111100",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0111111100",
		"0111111100",
		"0111111000",
		"0110011100",
		"0110001100",
		"0110001100",
		"0110000110",
		"0110000110",
		"0110000110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--R}
		--{S
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0011111100",
		"0011111100",
		"0110000110",
		"0110000110",
		"0110000110",
		"0011000000",
		"0011000000",
		"0001111000",
		"0000001100",
		"0000001100",
		"0110000110",
		"0110000110",
		"0110000110",
		"0011111100",
		"0011111100",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--S}
		--{T
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0111111110",
		"0111111110",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--T}
		--{U
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0011111100",
		"0011111100",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--U}
		--{V
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0011001100",
		"0011001100",
		"0011001100",
		"0011001100",
		"0011001100",
		"0011001100",
		"0011001100",
		"0001111000",
		"0000110000",
		"0000110000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--V}
		--{W
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110110110",
		"0110110110",
		"0111001110",
		"0111001110",
		"0110000110",
		"0110000110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--W}
		--{X
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0110000110",
		"0110000110",
		"0110000110",
		"0011001100",
		"0011001100",
		"0011001100",
		"0000110000",
		"0000110000",
		"0000110000",
		"0011001100",
		"0011001100",
		"0011001100",
		"0110000110",
		"0110000110",
		"0110000110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--X}
		--{Y
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0110000110",
		"0110000110",
		"0011001100",
		"0011001100",
		"0011001100",
		"0001111000",
		"0001111000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--Y}
		--{Z
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0111111110",
		"0111111110",
		"0000000110",
		"0000000110",
		"0000000110",
		"0000001100",
		"0000011100",
		"0001111000",
		"0011100000",
		"0011000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0111111110",
		"0111111110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--Z}
		--{[
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0111111110",
		"0111111110",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0111111110",
		"0111111110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--[}
		--{\
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"1100000000",
		"1100000000",
		"1100000000",
		"0011000000",
		"0011000000",
		"0011000000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000001100",
		"0000001100",
		"0000001100",
		"0000000011",
		"0000000011",
		"0000000011",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--\}
		--{]
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0111111110",
		"0111111110",
		"0000000110",
		"0000000110",
		"0000000110",
		"0000000110",
		"0000000110",
		"0000000110",
		"0000000110",
		"0000000110",
		"0000000110",
		"0000000110",
		"0000000110",
		"0111111110",
		"0111111110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--]}
		--{^
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000110000",
		"0001111000",
		"0011001100",
		"0110000110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--^}
		--{_
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"1111111111",
		"1111111111",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--_}
		--{`
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		
		"0111100000",
		"0111100000",
		"0001100000",
		"0001100000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--`}
		--{a
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0001111100",
		"0011111110",
		"0000000110",
		"0011111110",
		"0111111110",
		"0110000110",
		"0110000110",
		"0111111110",
		"0011110110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--a}
		--{b
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0111111100",
		"0111111110",
		"0110000110",
		"0110000110",
		"0111111110",
		"0110111100",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--b}
		--{c
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0011111100",
		"0111111110",
		"0110000110",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000110",
		"0111111110",
		"0011111100",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--c}
		--{d
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000110",
		"0000000110",
		"0000000110",
		"0011111110",
		"0111111110",
		"0110000110",
		"0110000110",
		"0111111110",
		"0011110110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--d}
		--{e
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0011111100",
		"0111111110",
		"0110000110",
		"0110000110",
		"0111111110",
		"0111111110",
		"0110000000",
		"0110000110",
		"0011111100",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--e}
		--{f
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0001111110",
		"0011111110",
		"0011000000",
		"0111111110",
		"0111111110",
		"0011000000",
		"0011000000",
		"0011000000",
		"0011000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--f}
		--{g
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0011110110",
		"0111111110",
		"0110000110",
		"0111111110",
		"0011111110",
		"0000000110",
		"0110000110",
		"0111111110",
		"0011111100",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--g}
		--{h
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0111111100",
		"0111111110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--h}
		--{i
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000110000",
		"0000110000",
		"0000000000",
		"0000000000",
		"0001110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0001111000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--i}
		--{j
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000110",
		"0000000110",
		"0000000000",
		"0000001110",
		"0000000110",
		"0000000110",
		"0110000110",
		"0111111110",
		"0011111100",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--j}
		--{k
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0110000000",
		"0110000000",
		"0110000110",
		"0110000110",
		"0111111100",
		"0110110000",
		"0110011000",
		"0110001100",
		"0110000110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--k}
		--{l
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0001110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0001111000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--l}
		--{m
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0011001100",
		"0111111110",
		"0110110110",
		"0110110110",
		"0110110110",
		"0110110110",
		"0110110110",
		"0110110110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--m}
		--{n
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0110111100",
		"0111111110",
		"0111000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--n}
		--{o
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0011111100",
		"0111111110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0111111110",
		"0011111100",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--o}
		--{p
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0110111100",
		"0111111110",
		"0110000110",
		"0110000110",
		"0111111110",
		"0111111100",
		"0110000000",
		"0110000000",
		"0110000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--p}
		--{q
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0011110110",
		"0111111110",
		"0110000110",
		"0110000110",
		"0111111110",
		"0011110110",
		"0000000110",
		"0000000110",
		"0000000110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--q}
		--{r
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0110111100",
		"0111111110",
		"0110000110",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0110000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--r}
		--{s
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0011111100",
		"0111111110",
		"0110000110",
		"0110000000",
		"0011111100",
		"0000000110",
		"0110000110",
		"0111111110",
		"0011111100",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--s}
		--{t
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0011000000",
		"0111111110",
		"0111111110",
		"0011000000",
		"0011000000",
		"0011000000",
		"0011000110",
		"0011111110",
		"0001111100",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--t}
		--{u
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0111111110",
		"0011110110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--u}
		--{v
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0011001100",
		"0011001100",
		"0001111000",
		"0000110000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--v}
		--{w
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110000110",
		"0110110110",
		"0110110110",
		"0011001100",
		"0011001100",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--w}
		--{x
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0110000110",
		"0110000110",
		"0011001100",
		"0001111000",
		"0000110000",
		"0001111000",
		"0011001100",
		"0110000110",
		"0110000110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--x}
		--{y
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0110000110",
		"0110000110",
		"0110000110",
		"0111111110",
		"0011111110",
		"0000000110",
		"0110000110",
		"0111111110",
		"0011111100",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--y}
		--{z
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0111111110",
		"0111111110",
		"0000000110",
		"0000011100",
		"0001111000",
		"0011100000",
		"0110000000",
		"0111111110",
		"0111111110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--z}
		--{{
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0001111110",
		"0011111110",
		"0011000000",
		"0011000000",
		"0011000000",
		"0011000000",
		"0011000000",
		"0110000000",
		"0011000000",
		"0011000000",
		"0011000000",
		"0011000000",
		"0011000000",
		"0011111110",
		"0001111110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--{}
		--{|
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--|}
		--{}
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0111111000",
		"0111111100",
		"0000001100",
		"0000001100",
		"0000001100",
		"0000001100",
		"0000001100",
		"0000000110",
		"0000001100",
		"0000001100",
		"0000001100",
		"0000001100",
		"0000001100",
		"0111111100",
		"0111111000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--}}
		--{~
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0111100000",
		"1100110011",
		"0000011110",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--~}
		--{DEL
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--DEL}
		-- skipping some of the extended ascii codes
		-- only including a few drawing chars
		-- sigle line box chars, and fill chars
		--{ bottom right corner (128)
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"1111110000",
		"1111110000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--}
		--{ top right corner (129)
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"1111110000",
		"1111110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		--}
		--{ top left corner (130)
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000111111",
		"0000111111",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		--}
		--{ bottom left corner (131)
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000111111",
		"0000111111",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		--}
		--{ cross (132)
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"1111111111",
		"1111111111",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		--}
		--{ horizontal line (133)
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"1111111111",
		"1111111111",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--}
		--{ right tee (134)
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000111111",
		"0000111111",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		--}
		--{ left tee (135)
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"1111110000",
		"1111110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		--}
		--{ up tee (136)
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"1111111111",
		"1111111111",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--}
		--{ down tee (137)
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"1111111111",
		"1111111111",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		--}
		--{ vertical line (138)
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		"0000110000",
		--}
		--{ quarter fill (139)
		"1100110011",
		"1100110011",
		"0011001100",
		"0011001100",
		"1100110011",
		"1100110011",
		"0011001100",
		"0011001100",
		"1100110011",
		"1100110011",
		"0011001100",
		"0011001100",
		"1100110011",
		"1100110011",
		"0011001100",
		"0011001100",
		"1100110011",
		"1100110011",
		"0011001100",
		"0011001100",
		"1100110011",
		"1100110011",
		"0011001100",
		"0011001100",
		"0011001100",
		--}
		--{ half fill (140)
		"1010101010",
		"0101010101",
		"1010101010",
		"0101010101",
		"1010101010",
		"0101010101",
		"1010101010",
		"0101010101",
		"1010101010",
		"0101010101",
		"1010101010",
		"0101010101",
		"1010101010",
		"0101010101",
		"1010101010",
		"0101010101",
		"1010101010",
		"0101010101",
		"1010101010",
		"0101010101",
		"1010101010",
		"0101010101",
		"1010101010",
		"0101010101",
		"1010101010",
		--}
		--{ full block (141)
		"1111111111",
		"1111111111",
		"1111111111",
		"1111111111",
		"1111111111",
		"1111111111",
		"1111111111",
		"1111111111",
		"1111111111",
		"1111111111",
		"1111111111",
		"1111111111",
		"1111111111",
		"1111111111",
		"1111111111",
		"1111111111",
		"1111111111",
		"1111111111",
		"1111111111",
		"1111111111",
		"1111111111",
		"1111111111",
		"1111111111",
		"1111111111",
		"1111111111",
		--}
		--{ cursor (142)
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"1111111111",
		"1111111111",
		"1111111111",
		"1111111111",
		"1111111111",
		"1111111111",
		"1111111111",
		"1111111111",
		"1111111111",
		"1111111111",
		"1111111111",
		"1111111111",
		"1111111111",
		"1111111111",
		"1111111111",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		"0000000000",
		--}
		others => "0000000000"
	);

end architecture a0;